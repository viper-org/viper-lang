struct abc {
    test: i32[3];
    foo: i32;
}